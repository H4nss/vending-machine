LIBRARY ieee;
use ieee.std_logic_1164.all;

package resource_holder_pkg is

    component resource_holder
        port()

end package resource_holder_pkg;

